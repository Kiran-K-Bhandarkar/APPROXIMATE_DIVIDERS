LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL; 

ENTITY DIVIDER_TB IS
END ENTITY DIVIDER_TB;

ARCHITECTURE TEST OF DIVIDER_TB IS
-----------------------------------------------------------------------------
  -- TESTBENCH INTERNAL SIGNALS
-----------------------------------------------------------------------------
CONSTANT DT_WIDTH: INTEGER := 16;
CONSTANT TFT_WIDTH: INTEGER := 8;
CONSTANT CLK_PERIOD: TIME := 5 NS; 
FILE FILE_VECTORS : TEXT;
FILE FILE_RESULTS : TEXT;
SIGNAL CLK, RST: STD_LOGIC;
SIGNAL IN1: STD_LOGIC_VECTOR(DT_WIDTH-1 DOWNTO 0);
SIGNAL IN2, QNT, RE: STD_LOGIC_VECTOR((DT_WIDTH/2)-1 DOWNTO 0);

BEGIN
  UUT: ENTITY WORK.DIVIDER_TM
    GENERIC MAP (DIVIDER_WIDTH => DT_WIDTH, TUNING_FACTOR => TFT_WIDTH)
	PORT MAP (CLK => CLK, RST => RST, IN1 => IN1, IN2 => IN2, QNT => QNT, RE => RE);
  
  CLK_PROCESS: PROCESS
   BEGIN
	CLK <= '1';
	WAIT FOR CLK_PERIOD/2;
	CLK <= '0';
	WAIT FOR CLK_PERIOD/2;
   END PROCESS CLK_PROCESS;	
   
  TEST_PROCESS: PROCESS
    VARIABLE V_ILINE     : LINE;
    VARIABLE V_OLINE     : LINE;
	VARIABLE V_SPACE     : CHARACTER;
    VARIABLE V_DIVIDEND  : INTEGER;
    VARIABLE V_DIVISOR   : INTEGER;
	
   BEGIN
    FILE_OPEN(FILE_VECTORS, "DIVIDER_INPUT.TXT", READ_MODE);
	FILE_OPEN(FILE_RESULTS, "DIVIDER_OUTPUT.TXT", WRITE_MODE);
	
	RST <= '1';
	WAIT FOR CLK_PERIOD;
	RST <= '0';
	WAIT FOR CLK_PERIOD;
	
   WHILE NOT ENDFILE(FILE_VECTORS) LOOP
      READLINE(FILE_VECTORS, V_ILINE);
      READ(V_ILINE, V_DIVIDEND);
      READ(V_ILINE, V_SPACE);          
      READ(V_ILINE, V_DIVISOR);
 
      IN1 <= STD_LOGIC_VECTOR(TO_UNSIGNED(V_DIVIDEND, IN1'LENGTH));
      IN2 <= STD_LOGIC_VECTOR(TO_UNSIGNED(V_DIVISOR, IN2'LENGTH));
 
      WAIT FOR CLK_PERIOD/2;
	  
      WRITE(V_OLINE, TO_INTEGER(UNSIGNED(QNT)));
	  WRITE(V_OLINE, V_SPACE);
      WRITE(V_OLINE, TO_INTEGER(UNSIGNED(RE)));
	  WRITELINE(FILE_RESULTS, V_OLINE);
	  
	  WAIT FOR CLK_PERIOD/2;
   END LOOP;
	  FILE_CLOSE(FILE_VECTORS);
	  FILE_CLOSE(FILE_RESULTS);
      WAIT;
   END PROCESS TEST_PROCESS;
END ARCHITECTURE TEST;