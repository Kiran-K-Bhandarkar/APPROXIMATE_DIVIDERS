LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DIVIDER_TM IS
GENERIC
(
	DIVIDER_WIDTH: INTEGER := 16;
	TUNING_FACTOR: INTEGER := 8
);
PORT
(
	CLK, RST: IN STD_LOGIC;
	IN1: IN STD_LOGIC_VECTOR(DIVIDER_WIDTH-1 DOWNTO 0);
	IN2: IN STD_LOGIC_VECTOR((DIVIDER_WIDTH/2)-1 DOWNTO 0);
	QNT: OUT STD_LOGIC_VECTOR((DIVIDER_WIDTH/2)-1 DOWNTO 0);
	RE: OUT STD_LOGIC_VECTOR((DIVIDER_WIDTH/2)-1 DOWNTO 0)
);
END ENTITY DIVIDER_TM;

ARCHITECTURE STRUCT OF DIVIDER_TM IS
CONSTANT D_WIDTH: INTEGER := DIVIDER_WIDTH;
CONSTANT T_FACTOR: INTEGER := TUNING_FACTOR;
SIGNAL Z_TEMP: STD_LOGIC_VECTOR(D_WIDTH-1 DOWNTO 0);
SIGNAL D_TEMP: STD_LOGIC_VECTOR((D_WIDTH/2)-1 DOWNTO 0);
SIGNAL Q_TEMP: STD_LOGIC_VECTOR((D_WIDTH/2)-1 DOWNTO 0);
SIGNAL S_TEMP: STD_LOGIC_VECTOR((D_WIDTH/2)-1 DOWNTO 0);

BEGIN
  REG_DIVID: ENTITY WORK.REG 
	  GENERIC MAP (INPUT_WIDTH => D_WIDTH)
	  PORT MAP
		(
		  CLK => CLK,
		  RST => RST,
		  INPUT => IN1,
		  OUTPUT => Z_TEMP
		);
	
	REG_DIVIS: ENTITY WORK.REG
	  GENERIC MAP (INPUT_WIDTH => D_WIDTH/2)
	  PORT MAP
		(
		  CLK => CLK,
		  RST => RST,
		  INPUT => IN2,
		  OUTPUT => D_TEMP
		);
	
	REG_QNT: ENTITY WORK.REG 
	  GENERIC MAP (INPUT_WIDTH => D_WIDTH/2)
	  PORT MAP
		(
		  CLK => CLK,
		  RST => RST,
		  INPUT => Q_TEMP,
		  OUTPUT => QNT
		);
		
	REG_REM: ENTITY WORK.REG 
	  GENERIC MAP (INPUT_WIDTH => D_WIDTH/2)
	  PORT MAP
		(
		  CLK => CLK,
		  RST => RST,
		  INPUT => S_TEMP,
		  OUTPUT => RE
		);
	
	DIV: ENTITY WORK.DIVIDER
	  GENERIC MAP (DIVIDER_WIDTH => D_WIDTH, TUNING_FACTOR => T_FACTOR)
	  PORT MAP
	    (
	     Z => Z_TEMP,
		  D => D_TEMP,
		  Q => Q_TEMP,
		  S => S_TEMP
	    );
END ARCHITECTURE STRUCT;
	  
